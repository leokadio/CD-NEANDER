library verilog;
use verilog.vl_types.all;
entity ldm_neander_vlg_vec_tst is
end ldm_neander_vlg_vec_tst;
