library verilog;
use verilog.vl_types.all;
entity ldm_controle_neander_vlg_vec_tst is
end ldm_controle_neander_vlg_vec_tst;
