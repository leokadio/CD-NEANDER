library verilog;
use verilog.vl_types.all;
entity ldm_fsm_tp8_vlg_vec_tst is
end ldm_fsm_tp8_vlg_vec_tst;
