library verilog;
use verilog.vl_types.all;
entity ldm_counter_8bits_vlg_vec_tst is
end ldm_counter_8bits_vlg_vec_tst;
